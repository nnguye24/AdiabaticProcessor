module CU_tb();





endmodule