module sram_bank_tb();


initial begin
    $dumpfile("sram_bank.vcd");
    $dumpvars(0, bank_tb);
end
endmodule